module ripple_carry_adder_4bit(
    input  logic [3:0] A,
    input  logic [3:0] B,
    input  logic Cin,
    output logic [3:0] S,
    output logic Cout
);
endmodule